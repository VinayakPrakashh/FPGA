`timescale 1ns / 1ps
module top(
clk,rst
    );
//inputs
input clk,rst;



//wire

endmodule
